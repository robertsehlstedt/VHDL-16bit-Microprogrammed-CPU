-- umem.vhd
-- This file implements the micro memory of the computer.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity umem is
  port(
    adr :       in std_logic_vector(7 downto 0)         := (others => '0');
    data :      out std_logic_vector(29 downto 0)       := (others => '0')
    );
end umem;

architecture behaviour of umem is
  type u_mem_t is array (0 to 255) of std_logic_vector(29 downto 0);

  -- MICRO MEMORY
  constant u_mem_c : u_mem_t :=
    -- _ALU__TB___FB__R__SP_PC_I_SEQ___uAddr
    (b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_1_0000_00000000",  -- 00, IR=PM(PC)
     b"0000_0000_0000_00_00_1_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0010_00000000",  -- uPC=K2
     
     b"1101_0110_0001_11_00_1_0_0001_00000000",  -- 04, IMMEDIATE AR=PM
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",  
     b"0000_0000_0000_00_00_0_0_0000_00000000",  

     b"0000_0110_0010_10_00_0_0_0000_00000000",  -- 08, Direct, ADR=IR(8 bits), PC++
     b"1101_1001_0001_00_00_0_0_0001_00000000",  -- AR=DM(ADR), uPC=K1
     b"0000_0110_0010_10_00_0_0_0000_00000000",  -- Indirect, ADR=IR(8 bits), PC++
     b"0000_1001_0010_00_00_0_0_0000_00000000",  -- ADR=DM(ADR)

     b"1101_1001_0001_00_00_0_0_0001_00000000",  -- 0C, AR=DM(ADR), uPC=K1
     b"0000_0011_0101_00_00_0_0_0011_00000000",  -- ((JMP))
     b"0000_0011_0111_00_00_0_0_0011_00000000",  -- ((LD))
     b"0000_0111_1000_01_00_0_0_0000_00000000",  -- ((CPY))

     b"0000_1000_0111_00_00_0_0_0011_00000000",  -- 10
     b"0000_0011_1001_00_00_0_0_0011_00000000",  -- ((STI))
     b"0000_0111_1001_00_00_0_0_0011_00000000",  -- ((ST))
     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- ((CMP))

     b"0010_0111_0001_00_00_0_0_0011_00000000",  -- 14
     b"0000_0111_1000_00_00_0_0_0000_00000000",  -- ((SWP))
     b"1101_0111_0001_01_00_0_0_0000_00000000",
     b"0000_0011_0111_00_00_0_0_0000_00000000",

     b"0000_1000_0111_01_00_0_0_0011_00000000",  -- 18
     b"0000_0100_0010_00_01_0_0_0000_00000000",  -- ((CALL))
     b"0000_0101_1001_00_00_0_0_0000_00000000",
     b"0000_0011_0101_00_00_0_0_0011_00000000",

     b"0000_0000_0000_00_10_0_0_0000_00000000",  -- 1C ((RET))
     b"0000_0100_0010_00_00_0_0_0000_00000000",
     b"0000_1001_0101_00_00_0_0_0011_00000000",
     b"0000_0000_0000_00_00_0_0_1000_00001101",  -- ((BEQ))

     b"0000_0000_0000_00_00_0_0_0011_00000000",  -- 20
     b"0000_0000_0000_00_00_0_0_1000_00000000",  -- ((BNE))
     b"0000_0000_0000_00_00_0_0_0100_00001101",
     b"0000_0000_0000_00_00_0_0_1010_00000000",  -- ((BCC))

     b"0000_0000_0000_00_00_0_0_0100_00001101",  -- 24
     b"0000_0000_0000_00_00_0_0_1010_00001101",  -- ((BCS))
     b"0000_0000_0000_00_00_0_0_0011_00000000",
     b"0000_0000_0000_00_00_0_0_1001_00001101",  -- ((BMI))

     b"0000_0000_0000_00_00_0_0_0011_00000000",  -- 28
     b"0000_0000_0000_00_00_0_0_1001_00000000",  -- ((BPL))
     b"0000_0000_0000_00_00_0_0_0100_00001101",
     b"0000_0000_0000_00_00_0_0_1011_00000000",  -- ((BVC))

     b"0000_0000_0000_00_00_0_0_0100_00001101",  -- 2C
     b"0000_0000_0000_00_00_0_0_1011_00001101",  -- ((BVS))
     b"0000_0000_0000_00_00_0_0_0011_00000000",
     b"1101_0111_0001_00_00_0_0_0000_00000000",  -- ((ADD))

     b"0001_0111_0001_01_00_0_0_0000_00000000",  -- 30
     b"0000_0011_0111_00_00_0_0_0011_00000000",
     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- ((SUB))
     b"0010_0111_0001_00_00_0_0_0000_00000000",

     b"0000_0011_0111_00_00_0_0_0011_00000000",  -- 34
     b"1101_0111_0001_00_00_0_0_0000_00000000",  -- ((AND))
     b"0111_0111_0001_01_00_0_0_0000_00000000",
     b"0000_0011_0111_00_00_0_0_0011_00000000",

     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- 38 ((OR))
     b"1000_0111_0001_00_00_0_0_0000_00000000",
     b"0000_0011_0111_00_00_0_0_0011_00000000",
     b"1001_0111_0001_00_00_0_0_0000_00000000",  -- ((LSL))

     b"0000_0011_0111_00_00_0_0_0011_00000000",  -- 3C
     b"1010_0111_0001_00_00_0_0_0000_00000000",  -- ((LSR))
     b"0000_0011_0111_00_00_0_0_0011_00000000",
     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- ((MUL))

     b"0011_0111_0001_00_00_0_0_0000_00000000",  -- 40
     b"0000_0011_0111_00_00_0_0_0011_00000000",
     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- ((MULS))
     b"0100_0111_0001_00_00_0_0_0000_00000000",

     b"0000_0011_0111_00_00_0_0_0011_00000000",  -- 44
     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- ((DIV))
     b"0101_0111_0001_00_00_0_0_0000_00000000",
     b"0000_0011_0111_00_00_0_0_0011_00000000",

     b"1101_0111_0001_01_00_0_0_0000_00000000",  -- 48 ((DIVS))
     b"0110_0111_0001_00_00_0_0_0000_00000000",
     b"0000_0011_0111_00_00_0_0_0011_00000000",
     b"1100_0111_0001_00_00_0_0_0000_00000000",  -- ((COM))

     b"0000_0011_0111_00_00_0_0_0011_00000000",  -- 4C
     b"0000_0111_1010_00_00_0_0_0000_00000000",  -- ((DRW))
     b"0000_0111_1011_01_00_0_0_0000_00000000",
     b"0000_0011_1100_00_00_0_0_0011_00000000",

     b"0000_0011_1100_00_00_0_0_0011_00000000",  -- 50 ((FWDB))
     b"0000_0011_1101_00_00_0_0_0000_00000000",  -- ((KBD))
     b"1101_1110_0001_00_00_0_0_0011_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",  -- 54
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",  -- 58
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",  -- 5C
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",  -- 60
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",  -- 64
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",  -- 68
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 6C
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 70
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 74
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 78
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 7C
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 80
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 84
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 88
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 8C
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 80
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 94
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 98
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- 9C
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- A0
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- A4
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- A8
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- AC
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- B0
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- B4
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- B8
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- BC
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- C0
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- C4
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- C8
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- CC
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- D0
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- D4
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- D8
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- DC
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- E0
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- E4
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- E8
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- EC
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- F0
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- F4
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- F8
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",

     b"0000_0000_0000_00_00_0_0_0000_00000000",       -- FC
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0000_00000000",
     b"0000_0000_0000_00_00_0_0_0001_00000000"        -- (When no mode
                                                      -- necessary,uPC=K1, PC++)
     );

  signal u_mem : u_mem_t := u_mem_c;

  begin
    data <= u_mem(to_integer(unsigned(adr)));
end architecture behaviour;
